LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DATA_PATH IS 
PORT 
(
CARGA_DATA_REGISTRO :  STD_LOGIC_VECTOR (7 DOWNTO 0);
 SALIDA_B : BUFFER STD_LOGIC_VECTOR (3 DOWNTO 0);
Z_NOR, A_SALIDA : BUFFER STD_LOGIC;
 L, E, LB, EB : IN STD_LOGIC;
CLOCK_PULSADOR : IN STD_LOGIC
);
END DATA_PATH;

ARCHITECTURE ARQUI OF DATA_PATH IS
 

COMPONENT CONTADOR_CON_DATO IS 
------------------------------
--DECLARAREMOS LAS VARIABLES
GENERIC(VARIABLE1 : INTEGER := 4);
PORT 
(
RELOJ_DE_ENTRADA, ENABLE: IN STD_LOGIC;
CARGA_PARALELA : IN STD_LOGIC;
CARGA_PARALELA_DATO : IN STD_LOGIC_VECTOR (VARIABLE1 - 1 DOWNTO 0); 
CONTADOR_SALIDA : BUFFER STD_LOGIC_VECTOR (VARIABLE1 - 1 DOWNTO 0)
);
END COMPONENT;

-----------------------------------

COMPONENT shiftregRight_syncLoad IS

GENERIC(		N  : INTEGER:= 8	);

PORT
 (
	clk								:  IN  STD_LOGIC;									-- RELOJ DE SHIFT REGISTER
	DataIn							:  IN  STD_LOGIC;									-- SERIAL DATA
   enableShift, enableLoad 	: 	IN  STD_LOGIC;									--	ENTRADAS SHIFT, ENABLE SYNC LOAD RESPECTIVELY
	dataLoad							:  IN  STD_LOGIC_VECTOR(N-1 DOWNTO 0);		-- LOADING DATA
	q		  							: 	OUT std_logic_VECTOR(N-1 DOWNTO 0)
); 	-- PARALLEL OUTPUTS SHIFT REGISTER

END COMPONENT;

----------------------------------

 SIGNAL SALIDA_Q : STD_LOGIC_VECTOR (7 DOWNTO 0);
 SIGNAL CARGA_CONTADOR: STD_LOGIC_VECTOR ( 3 DOWNTO 0) := "0000";
 
BEGIN

REGISTRO: shiftregRight_syncLoad PORT MAP ( dataLoad => CARGA_DATA_REGISTRO, DataIn => '0', clk => CLOCK_PULSADOR, q => SALIDA_Q, enableShift => E, enableLoad => L );

A_SALIDA <= SALIDA_Q(0);

Z_NOR <= NOT(SALIDA_Q(7) OR SALIDA_Q(6) OR SALIDA_Q(5) OR SALIDA_Q(4) OR SALIDA_Q(3) OR SALIDA_Q(2) OR SALIDA_Q(1) OR SALIDA_Q(0));

COUNTER: CONTADOR_CON_DATO PORT MAP ( CARGA_PARALELA_DATO => CARGA_CONTADOR, RELOJ_DE_ENTRADA => CLOCK_PULSADOR, ENABLE => EB, CARGA_PARALELA => LB, CONTADOR_SALIDA => SALIDA_B );

END ARQUI;