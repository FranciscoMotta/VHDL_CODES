LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY divisor_50_to_1k IS 
PORT 
( 
SALIDA: BUFFER STD_LOGIC;
CLK_IN: IN STD_LOGIC
);
END divisor_50_to_1k;


ARCHITECTURE DIVISOR_DE_FREQ OF divisor_50_to_1k IS
CONSTANT TOP: STD_LOGIC_VECTOR (27 DOWNTO 0) := x"0001387"; 
SIGNAL CONTADOR : STD_LOGIC_VECTOR (27 DOWNTO 0) := x"0000000";
SIGNAL CLK_OUT: STD_LOGIC;
BEGIN 
PROCESS (CLK_IN)
BEGIN
	IF(CLK_IN'EVENT AND CLK_IN ='1') THEN

	--DISEÃ‘O DEL CONTADOR
	 
	  IF (CONTADOR = TOP) THEN 
	  CONTADOR <= x"0000000";
	  ELSE 
		CONTADOR <= CONTADOR + x"0000001";
	  END IF;
	  
	--DISEÃ‘O DEL COMPARADOR

		IF (CONTADOR = TOP) THEN 
			SALIDA <= '1';
		ELSE 
			SALIDA <= '0';
		END IF;	
	END IF;
END PROCESS;


END DIVISOR_DE_FREQ;