LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALGORITMOS IS
PORT
(
CARGA_CONTADOR : INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
DATA : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
SALIDA_B : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
);
END ALGORITMOS;

ARCHITECTURE ARQUI OF ALGORITMOS IS 

--------------------------------------

----------------COMPONENTES--------------

COMPONENT divisor_50_to_1k IS 
PORT 
( 
SALIDA: BUFFER STD_LOGIC;
CLK_IN: IN STD_LOGIC
);
END COMPONENT;


--------------------------------

---------DECLARACION DE SEÑALES



BEGIN 

END ARQUI;